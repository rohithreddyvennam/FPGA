module qpsktest(
	input clk,
	input [7:0] x_in,
	output [3:0] y_out
);

  reg [3:0] temp;

  initial begin
	temp <= 8'd0;
  end
  
  assign y_out = ~temp;

  always@(posedge clk) begin
	temp[0] <= x_in[0];
	temp[1] <= x_in[2];
	temp[2] <= x_in[4];
	temp[3] <= x_in[6];
  end

endmodule
	
